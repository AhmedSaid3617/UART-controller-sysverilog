module uart_controller ();

    

endmodule

