interface uart_rx_if;
    
endinterface

module uart_rx ();
    
endmodule